interface and_if();

	logic p,r;
	logic r;
	modport  dut_mp(input p,input q,output r);
	modport  tb_mp(input p,input  q,output r);
	

endinterface
