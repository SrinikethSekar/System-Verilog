module design(and_if inst);

	assign inst.dut_mp.r=inst.dut_mp.p & inst.dut_mp.q;

endmodule
