module and_i(and_if inst);

	assign inst.ans=inst.a&inst.b;


endmodule
