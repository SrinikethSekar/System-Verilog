interface and_if;

	logic a;
	logic b;
	logic ans;



endinterface
