module r_case;

  initial begin   

    $display("INDIAN CRICKET");
    $display("ALAPARAI");
    
    for (int i = 0; i < 6; i++) begin

      randcase

        0: $display("\t \n Thala sons"); 
        1: $display("\t \n Virat Veriyans"); 
        2: $display("\t \n Rohit Fans muttu"); 
        3: $display("\t \n Gambir fans credit");
      
      endcase

    end

  end

endmodule


// INDIAN CRICKET
// ALAPARAI
   
//  Rohit Fans muttu
   
//  Gambir fans credit
   
//  Virat Veriyans
   
//  Gambir fans credit
   
//  Gambir fans credit
   
//  Gambir fans credit
